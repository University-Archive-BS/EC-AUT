** Profile: "SCHEMATIC1-pish_gozaresh"  [ D:\DOCUMENTS\POLYTECHNIC\TERM 3\ELECTRICAL CIRCUITS LAB\AZ4\AZ4 Q4\pish_gozaresh-SCHEMATIC1-pish_gozaresh.sim ] 

** Creating circuit file "pish_gozaresh-SCHEMATIC1-pish_gozaresh.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 .1s 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pish_gozaresh-SCHEMATIC1.net" 


.END
