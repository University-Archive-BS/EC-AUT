** Profile: "SCHEMATIC1-AZ4"  [ d:\documents\polytechnic\term 3\electrical circuits lab\az4 q1s2\az4-schematic1-az4.sim ] 

** Creating circuit file "az4-schematic1-az4.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V1 0 2V 0.1 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\az4-SCHEMATIC1.net" 


.END
