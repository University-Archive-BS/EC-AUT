** Profile: "SCHEMATIC1-AZ4Q1S1"  [ D:\DOCUMENTS\POLYTECHNIC\TERM 3\Electrical Circuits Lab\AZ4 Q1S1\az4q1s1-SCHEMATIC1-AZ4Q1S1.sim ] 

** Creating circuit file "az4q1s1-SCHEMATIC1-AZ4Q1S1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\az4q1s1-SCHEMATIC1.net" 


.END
