** Profile: "SCHEMATIC1-az10"  [ D:\DOCUMENTS\POLYTECHNIC\TERM 3\ELECTRICAL CIRCUITS LAB\AZ9\pish_gozaresh-SCHEMATIC1-az10.sim ] 

** Creating circuit file "pish_gozaresh-SCHEMATIC1-az10.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC LIN 200 100 1000
.OP
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pish_gozaresh-SCHEMATIC1.net" 


.END
