** Profile: "SCHEMATIC1-pishpish"  [ D:\DOCUMENTS\POLYTECHNIC\TERM 3\ELECTRICAL CIRCUITS LAB\AZ4\AZ4 Q4\pishgozaresh-SCHEMATIC1-pishpish.sim ] 

** Creating circuit file "pishgozaresh-SCHEMATIC1-pishpish.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 .1s 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pishgozaresh-SCHEMATIC1.net" 


.END
